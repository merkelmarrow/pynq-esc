`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: N/A
// Engineer: Marco Blackwell
// 
// Create Date: 16.08.2025 17:34:51
// Design Name: 
// Module Name: esc_mvp_top
// Project Name: PYNQ ESC
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module esc_mvp_top(
    input clk_125_in,
    input rst_n,
    output adc_mclk_out,
    output pwm_out
    );
    
    
endmodule
